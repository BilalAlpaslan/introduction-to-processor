module Ilk (A, B, C);
    output A, B, C;
    input X, Y, Z;
    wire W;
    and A, B, C;
endmodule